module MD (
    input   core_package:: md_op_e      opcode_i,
    input   logic [31:0]                operand_A_i,
    input   logic [31:0]                operand_B_i,
    output  logic [31:0]                result_o
);
    
endmodule