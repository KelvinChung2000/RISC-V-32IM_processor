module WB (
    ports
);
    
endmodule